Transient Analysis of CMOS Inverter
.Param supply = 5
VDD 3 0 supply
Mn 2 1 0 0 nmod w=10u l=1u
Mp 2 1 3 3 pmod w=20u l=1u
cload 2 0 1.5P
Vin 1 0 pulse(0 supply 8n 0 0 8n 16n)
.model NMOD NMOS VTO=1v kp=450u
.model PMOD PMOS VTO=1.2v kp=200u
.tran 1p 0.1u
.measure tran T_HL trig v(1) va1=2.5 rise=1 targ v(2) va1=2.5 fall=1
.measure tran T_LH trig v(1) va1=2.5 fall=1 targ v(2) va1=2.5 rise=1
.measure tran T_rise trig v(2) va1=0.5 rise=1 targ v(2) va1=4.5 rise=1
.measure tran T_fall trig v(2) va1=4.5 rise=1 targ v(2) va1=-0.5 fall=1
.control
run

set color0=white
set color1=blue
set color2=red
set color3=green

set xbrushwidth=2
plot v(2) v(2)+8
.endc
.end